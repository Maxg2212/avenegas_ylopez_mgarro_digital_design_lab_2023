module instruction_memory (
	input logic [31:0] a,
	output logic [31:0] rd
);

endmodule 